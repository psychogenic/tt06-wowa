magic
tech sky130A
magscale 1 2
timestamp 1712893257
<< pwell >>
rect -1083 -310 1083 310
<< nmos >>
rect -887 -100 -487 100
rect -429 -100 -29 100
rect 29 -100 429 100
rect 487 -100 887 100
<< ndiff >>
rect -945 88 -887 100
rect -945 -88 -933 88
rect -899 -88 -887 88
rect -945 -100 -887 -88
rect -487 88 -429 100
rect -487 -88 -475 88
rect -441 -88 -429 88
rect -487 -100 -429 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 429 88 487 100
rect 429 -88 441 88
rect 475 -88 487 88
rect 429 -100 487 -88
rect 887 88 945 100
rect 887 -88 899 88
rect 933 -88 945 88
rect 887 -100 945 -88
<< ndiffc >>
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
<< psubdiff >>
rect -1047 240 -951 274
rect 951 240 1047 274
rect -1047 178 -1013 240
rect 1013 178 1047 240
rect -1047 -240 -1013 -178
rect 1013 -240 1047 -178
rect -1047 -274 -951 -240
rect 951 -274 1047 -240
<< psubdiffcont >>
rect -951 240 951 274
rect -1047 -178 -1013 178
rect 1013 -178 1047 178
rect -951 -274 951 -240
<< poly >>
rect -887 172 -487 188
rect -887 138 -871 172
rect -503 138 -487 172
rect -887 100 -487 138
rect -429 172 -29 188
rect -429 138 -413 172
rect -45 138 -29 172
rect -429 100 -29 138
rect 29 172 429 188
rect 29 138 45 172
rect 413 138 429 172
rect 29 100 429 138
rect 487 172 887 188
rect 487 138 503 172
rect 871 138 887 172
rect 487 100 887 138
rect -887 -138 -487 -100
rect -887 -172 -871 -138
rect -503 -172 -487 -138
rect -887 -188 -487 -172
rect -429 -138 -29 -100
rect -429 -172 -413 -138
rect -45 -172 -29 -138
rect -429 -188 -29 -172
rect 29 -138 429 -100
rect 29 -172 45 -138
rect 413 -172 429 -138
rect 29 -188 429 -172
rect 487 -138 887 -100
rect 487 -172 503 -138
rect 871 -172 887 -138
rect 487 -188 887 -172
<< polycont >>
rect -871 138 -503 172
rect -413 138 -45 172
rect 45 138 413 172
rect 503 138 871 172
rect -871 -172 -503 -138
rect -413 -172 -45 -138
rect 45 -172 413 -138
rect 503 -172 871 -138
<< locali >>
rect -1047 240 -951 274
rect 951 240 1047 274
rect -1047 178 -1013 240
rect 1013 178 1047 240
rect -887 138 -871 172
rect -503 138 -487 172
rect -429 138 -413 172
rect -45 138 -29 172
rect 29 138 45 172
rect 413 138 429 172
rect 487 138 503 172
rect 871 138 887 172
rect -933 88 -899 104
rect -933 -104 -899 -88
rect -475 88 -441 104
rect -475 -104 -441 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 441 88 475 104
rect 441 -104 475 -88
rect 899 88 933 104
rect 899 -104 933 -88
rect -887 -172 -871 -138
rect -503 -172 -487 -138
rect -429 -172 -413 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 413 -172 429 -138
rect 487 -172 503 -138
rect 871 -172 887 -138
rect -1047 -240 -1013 -178
rect 1013 -240 1047 -178
rect -1047 -274 -951 -240
rect 951 -274 1047 -240
<< viali >>
rect -871 138 -503 172
rect -413 138 -45 172
rect 45 138 413 172
rect 503 138 871 172
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
rect -871 -172 -503 -138
rect -413 -172 -45 -138
rect 45 -172 413 -138
rect 503 -172 871 -138
<< metal1 >>
rect -883 172 -491 178
rect -883 138 -871 172
rect -503 138 -491 172
rect -883 132 -491 138
rect -425 172 -33 178
rect -425 138 -413 172
rect -45 138 -33 172
rect -425 132 -33 138
rect 33 172 425 178
rect 33 138 45 172
rect 413 138 425 172
rect 33 132 425 138
rect 491 172 883 178
rect 491 138 503 172
rect 871 138 883 172
rect 491 132 883 138
rect -939 88 -893 100
rect -939 -88 -933 88
rect -899 -88 -893 88
rect -939 -100 -893 -88
rect -481 88 -435 100
rect -481 -88 -475 88
rect -441 -88 -435 88
rect -481 -100 -435 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 435 88 481 100
rect 435 -88 441 88
rect 475 -88 481 88
rect 435 -100 481 -88
rect 893 88 939 100
rect 893 -88 899 88
rect 933 -88 939 88
rect 893 -100 939 -88
rect -883 -138 -491 -132
rect -883 -172 -871 -138
rect -503 -172 -491 -138
rect -883 -178 -491 -172
rect -425 -138 -33 -132
rect -425 -172 -413 -138
rect -45 -172 -33 -138
rect -425 -178 -33 -172
rect 33 -138 425 -132
rect 33 -172 45 -138
rect 413 -172 425 -138
rect 33 -178 425 -172
rect 491 -138 883 -132
rect 491 -172 503 -138
rect 871 -172 883 -138
rect 491 -178 883 -172
<< properties >>
string FIXED_BBOX -1030 -257 1030 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 2.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
