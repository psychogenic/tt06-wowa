magic
tech sky130A
magscale 1 2
timestamp 1713152285
<< error_s >>
rect -19013 -5000 -19000 -4800
rect -18985 -5000 -18972 -4772
<< metal1 >>
rect -18600 -200 -18400 0
rect -13400 -200 -13200 0
rect -11400 -200 -11200 0
rect -19200 -5000 -19000 -4800
rect -19200 -6000 -19000 -5800
rect -19200 -6400 -19000 -6200
rect -19200 -6800 -19000 -6600
rect -19200 -7200 -19000 -7000
rect -19200 -8000 -19000 -7800
use comparator_stefan  x1
timestamp 1713150544
transform 1 0 -28445 0 1 -10990
box 9445 5990 17870 10730
use analogswitch  x2
timestamp 1713149804
transform 1 0 -18620 0 1 -12120
box 5220 3520 7200 5620
use onehot2mux  x3
timestamp 1713137925
transform 1 0 -17650 0 1 -9780
box -550 1780 3445 3920
use sky130_fd_pr__cap_mim_m3_2_4HHTN9  XC1
timestamp 1713151418
transform 1 0 -8851 0 1 -4200
box -1349 -4800 1371 4800
<< labels >>
flabel metal1 -19200 -8000 -19000 -7800 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
flabel metal1 -19200 -5000 -19000 -4800 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
flabel metal1 -18600 -200 -18400 0 0 FreeSans 1280 0 0 0 VCC
port 0 nsew
flabel metal1 -13400 -200 -13200 0 0 FreeSans 1280 0 0 0 EN_N
port 6 nsew
flabel metal1 -11400 -200 -11200 0 0 FreeSans 1280 0 0 0 RESULT
port 5 nsew
flabel metal1 -19200 -7200 -19000 -7000 0 FreeSans 1280 0 0 0 THRESHV
port 3 nsew
flabel metal1 -19200 -6800 -19000 -6600 0 FreeSans 1280 0 0 0 INPUT
port 2 nsew
flabel metal1 -19200 -6400 -19000 -6200 0 FreeSans 1280 0 0 0 CALIB
port 4 nsew
flabel metal1 -19200 -6000 -19000 -5800 0 FreeSans 1280 0 0 0 VCC
port 0 nsew
<< end >>
