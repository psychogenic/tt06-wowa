* NGSPICE file created from wowa_analog.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_GGMWVD w_n996_n319# a_n800_n197# a_800_n100# a_n858_n100#
X0 a_800_n100# a_n800_n197# a_n858_n100# w_n996_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
**devattr s=11600,516 d=11600,516
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_3VR9VM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
**devattr s=11600,516 d=11600,516
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_FMMQLY a_100_n50# a_n100_n138# a_n260_n224# a_n158_n50#
X0 a_100_n50# a_n100_n138# a_n158_n50# a_n260_n224# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
**devattr s=5800,316 d=5800,316
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_FMHZDY a_n800_n138# a_n960_n224# a_n858_n50# a_800_n50#
X0 a_800_n50# a_n800_n138# a_n858_n50# a_n960_n224# sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
**devattr s=5800,316 d=5800,316
.ends

.subckt sky130_fd_pr__pfet_01v8_GGY9VD a_800_n200# a_n858_n200# w_n996_n419# a_n800_n297#
X0 a_800_n200# a_n800_n297# a_n858_n200# w_n996_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=8
**devattr s=23200,916 d=23200,916
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_GWPMZG a_n200_n897# a_200_n800# w_n396_n1019#
+ a_n258_n800#
X0 a_200_n800# a_n200_n897# a_n258_n800# w_n396_n1019# sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=2
**devattr s=92800,3316 d=92800,3316
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_FMZK9W a_400_n200# a_n458_n200# a_n400_n288# a_n560_n374#
X0 a_400_n200# a_n400_n288# a_n458_n200# a_n560_n374# sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=4
**devattr s=23200,916 d=23200,916
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD w_n596_n619# a_n400_n497# a_400_n400# a_n458_n400#
X0 a_400_n400# a_n400_n497# a_n458_n400# w_n596_n619# sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=4
**devattr s=46400,1716 d=46400,1716
.ends

.subckt sky130_fd_pr__pfet_01v8_UGSVTG a_15_n500# w_n211_n719# a_n33_n597# a_n73_n500#
X0 a_15_n500# a_n33_n597# a_n73_n500# w_n211_n719# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=0.15
**devattr s=58000,2116 d=58000,2116
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
.ends

.subckt comparator_stefan PLUS MINUS VCC VSS EN_N ADJ DIFFOUT
XXM12 VCC EN_N VCC p2p sky130_fd_pr__pfet_01v8_GGMWVD
XXM13 VCC ADJ G1 p2p sky130_fd_pr__pfet_01v8_lvt_3VR9VM
XXM14 G1 ADJ VSS n2n sky130_fd_pr__nfet_01v8_lvt_FMMQLY
XXM15 VCC VSS VSS n2n sky130_fd_pr__nfet_01v8_lvt_FMHZDY
XXM1 inhigh VCC VCC EN_N sky130_fd_pr__pfet_01v8_GGY9VD
XXM2 MINUS inhigh VCC G1 sky130_fd_pr__pfet_01v8_lvt_GWPMZG
XXM3 PLUS G2 VCC inhigh sky130_fd_pr__pfet_01v8_lvt_GWPMZG
XXM4 G2 VSS G2 VSS sky130_fd_pr__nfet_01v8_lvt_FMZK9W
XXM5 VSS G1 G1 VSS sky130_fd_pr__nfet_01v8_lvt_FMZK9W
XXM6 pg2g VSS G1 VSS sky130_fd_pr__nfet_01v8_lvt_FMZK9W
XXM7 VCC pg2g pg2g mirhigh sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD
XXM8 VCC pg2g mirhigh DIFFOUT sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD
XXM9 VCC VCC EN_N mirhigh sky130_fd_pr__pfet_01v8_UGSVTG
XXM10 VSS DIFFOUT G2 VSS sky130_fd_pr__nfet_01v8_lvt_FMZK9W
XXM11 DIFFOUT EN_N VSS VSS sky130_fd_pr__nfet_01v8_648S5X
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_4QFWD3 a_n93_n200# a_n35_n297# a_35_n200# w_n231_n419#
X0 a_35_n200# a_n35_n297# a_n93_n200# w_n231_n419# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.35
**devattr s=23200,916 d=23200,916
.ends

.subckt lvtnot a y VCCPIN VSUBS
XXM1 VSUBS a y VSUBS sky130_fd_pr__nfet_01v8_lvt_648S5X
XXM2 VCCPIN a y VCCPIN sky130_fd_pr__pfet_01v8_lvt_4QFWD3
.ends

.subckt sky130_fd_pr__nfet_01v8_Q7AWK3 a_n180_n374# a_20_n200# a_n78_n200# a_n33_n288#
X0 a_20_n200# a_n33_n288# a_n78_n200# a_n180_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
**devattr s=23200,916 d=23200,916
.ends

.subckt sky130_fd_pr__pfet_01v8_SKB8XJ w_n216_n419# a_n33_n297# a_20_n200# a_n78_n200#
X0 a_20_n200# a_n33_n297# a_n78_n200# w_n216_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
**devattr s=23200,916 d=23200,916
.ends

.subckt passgate A Z GP GN VCCBPIN VSUBS
XXM1 VSUBS Z A GN sky130_fd_pr__nfet_01v8_Q7AWK3
XXM2 VCCBPIN GP A Z sky130_fd_pr__pfet_01v8_SKB8XJ
.ends

.subckt analogswitch EN IN OUT VCC VSS
Xx1 EN x1/y VCC VSS lvtnot
Xx2 IN OUT x1/y EN VCC VSS passgate
.ends

.subckt onehot2mux SEL IN0 IN1 OUT VCC VSS
Xx1 SEL SEL_N VCC VSS lvtnot
Xx2 IN1 OUT SEL_N SEL VCC VSS passgate
Xx3 IN0 OUT SEL SEL_N VCC VSS passgate
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_4HHTN9 m3_n1186_n4520# c1_n1146_n4480#
X0 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X3 c1_n1146_n4480# m3_n1186_n4520# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt calibrated_comparator INPUT THRESHV RESULT EN_N CALIB VCC VSS
Xx1 x3/OUT THRESHV VCC VSS EN_N x2/OUT RESULT comparator_stefan
Xx2 CALIB RESULT x2/OUT VCC VSS analogswitch
Xx3 CALIB INPUT THRESHV x3/OUT VCC VSS onehot2mux
XXC1 VSS x2/OUT sky130_fd_pr__cap_mim_m3_1_4HHTN9
.ends

.subckt sky130_fd_pr__res_high_po_0p35_3KK54B a_n35_n4432# a_n35_4000# a_n165_n4562#
X0 a_n35_4000# a_n35_n4432# a_n165_n4562# sky130_fd_pr__res_high_po_0p35 l=40.16
.ends

.subckt sky130_fd_pr__res_high_po_0p35_QPS5FG a_n165_n2562# a_n35_n2432# a_n35_2000#
X0 a_n35_2000# a_n35_n2432# a_n165_n2562# sky130_fd_pr__res_high_po_0p35 l=20.16
.ends

.subckt r2r b0 b1 b2 b3 b4 b5 b6 b7 out VSUBS GND
XXR1 m1_n1840_11060# b0 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR10 VSUBS m1_n1040_2660# m1_n440_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR2 m1_n1040_2660# b1 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR11 VSUBS m1_160_2660# m1_n440_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR3 m1_n440_7180# b2 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR5 m1_760_7180# b4 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR12 VSUBS m1_160_2660# m1_760_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR4 m1_160_2660# b3 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR14 VSUBS m1_1360_2660# m1_1960_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR6 m1_1360_2660# b5 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR13 VSUBS m1_1360_2660# m1_760_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR15 VSUBS out m1_1960_7180# sky130_fd_pr__res_high_po_0p35_QPS5FG
XXR7 m1_1960_7180# b6 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR8 out b7 VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR16 GND m1_n1840_11060# VSUBS sky130_fd_pr__res_high_po_0p35_3KK54B
XXR9 VSUBS m1_n1040_2660# m1_n1840_11060# sky130_fd_pr__res_high_po_0p35_QPS5FG
.ends

.subckt wowa_analog b0 b1 b2 b3 b4 b5 b6 b7 EN_N CAL INPUT EXTTHRESH USEEXT VCC VSS
+ COMPOUT
Xx1 INPUT x3/OUT COMPOUT EN_N CAL VCC VSS calibrated_comparator
Xx2 b0 b1 b2 b3 b4 b5 b6 b7 x3/IN0 VSS VSS r2r
Xx3 USEEXT x3/IN0 EXTTHRESH x3/OUT VCC VSS onehot2mux
.ends

