magic
tech sky130A
magscale 1 2
timestamp 1713121489
<< nwell >>
rect -320 2020 -240 2120
<< pwell >>
rect -250 1670 -170 1690
rect -320 1580 -310 1590
rect -290 1580 -240 1590
rect -320 1570 -240 1580
rect -320 1500 -230 1570
<< viali >>
rect -380 2260 -30 2300
rect -380 1320 -40 1360
<< metal1 >>
rect -700 2300 300 2540
rect -700 2260 -380 2300
rect -30 2260 300 2300
rect -700 2240 300 2260
rect -250 2200 -240 2210
rect -700 2116 -500 2180
rect -260 2150 -240 2200
rect -180 2200 -170 2210
rect -180 2150 -160 2200
rect -700 2044 -516 2116
rect -444 2044 -438 2116
rect -700 1980 -500 2044
rect -340 2020 -240 2120
rect -180 2020 -80 2120
rect -340 1900 -280 2020
rect -250 1930 -240 1990
rect -180 1930 -170 1990
rect -140 1900 -80 2020
rect -700 1760 -280 1900
rect -150 1770 300 1900
rect -700 1730 -290 1760
rect -700 1700 -310 1730
rect -130 1720 300 1770
rect -700 1539 -500 1600
rect -340 1580 -310 1700
rect -110 1700 300 1720
rect -250 1680 -170 1690
rect -250 1620 -240 1680
rect -180 1620 -170 1680
rect -110 1580 -80 1700
rect -340 1570 -240 1580
rect -700 1462 -519 1539
rect -442 1462 -436 1539
rect -340 1500 -230 1570
rect -180 1500 -80 1580
rect -700 1400 -500 1462
rect -260 1400 -250 1470
rect -170 1400 -160 1470
rect -390 1360 -30 1370
rect -700 1320 -380 1360
rect -40 1320 300 1360
rect -700 1100 300 1320
<< via1 >>
rect -240 2150 -180 2210
rect -516 2044 -444 2116
rect -240 1930 -180 1990
rect -240 1620 -180 1680
rect -519 1462 -442 1539
rect -250 1400 -170 1470
<< metal2 >>
rect -240 2216 -180 2220
rect -246 2210 -174 2216
rect -246 2150 -240 2210
rect -180 2150 -174 2210
rect -516 2116 -444 2122
rect -246 2116 -174 2150
rect -444 2044 -174 2116
rect -516 2038 -444 2044
rect -246 1990 -174 2044
rect -246 1934 -240 1990
rect -180 1934 -174 1990
rect -240 1920 -180 1930
rect -250 1680 -170 1690
rect -250 1620 -240 1680
rect -180 1620 -170 1680
rect -250 1610 -170 1620
rect -519 1539 -442 1545
rect -249 1539 -172 1610
rect -442 1480 -172 1539
rect -442 1470 -170 1480
rect -442 1462 -250 1470
rect -519 1456 -442 1462
rect -250 1390 -170 1400
use sky130_fd_pr__nfet_01v8_L7T3GD  XM1
timestamp 1713118242
transform 1 0 -209 0 1 1542
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_M479BZ  XM2
timestamp 1713118242
transform 1 0 -209 0 1 2071
box -211 -261 211 261
<< labels >>
flabel metal1 -700 1400 -500 1600 0 FreeSans 1280 0 0 0 GN
port 3 nsew
flabel metal1 100 1700 300 1900 0 FreeSans 1280 0 0 0 Z
port 0 nsew
flabel metal1 -700 1700 -500 1900 0 FreeSans 1280 0 0 0 A
port 1 nsew
flabel metal1 -700 1980 -500 2180 0 FreeSans 1280 0 0 0 GP
port 2 nsew
flabel metal1 -300 2340 -100 2540 0 FreeSans 1280 0 0 0 VCCBPIN
port 4 nsew
flabel metal1 -400 1100 -200 1300 0 FreeSans 1280 0 0 0 VSSBPIN
port 5 nsew
<< end >>
