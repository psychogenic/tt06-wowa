magic
tech sky130A
magscale 1 2
timestamp 1712874608
<< metal1 >>
rect 28036 26414 28042 26474
rect 28102 26414 28108 26474
rect 28042 17758 28102 26414
rect 31356 21564 31362 21864
rect 31662 21564 31668 21864
rect 31362 17562 31662 21564
rect 28472 10790 28592 11332
rect 28466 10670 28472 10790
rect 28592 10670 28598 10790
rect 28476 10060 28482 10180
rect 28602 10060 28608 10180
rect 28482 9706 28602 10060
rect 29484 1882 29604 3776
rect 29688 1882 29808 1888
rect 29476 1762 29688 1882
rect 29688 1756 29808 1762
<< via1 >>
rect 28042 26414 28102 26474
rect 31362 21564 31662 21864
rect 28472 10670 28592 10790
rect 28482 10060 28602 10180
rect 29688 1762 29808 1882
<< metal2 >>
rect 31362 29587 31662 29592
rect 28042 29526 28102 29528
rect 28035 29470 28044 29526
rect 28100 29470 28109 29526
rect 28042 26474 28102 29470
rect 31358 29297 31367 29587
rect 31657 29297 31666 29587
rect 28042 26408 28102 26414
rect 31362 21864 31662 29297
rect 31362 21558 31662 21564
rect 26477 10790 26587 10794
rect 28472 10790 28592 10796
rect 26472 10785 28472 10790
rect 26472 10675 26477 10785
rect 26587 10675 28472 10785
rect 26472 10670 28472 10675
rect 26477 10666 26587 10670
rect 28472 10664 28592 10670
rect 28482 10180 28602 10186
rect 26896 10060 28482 10180
rect 26896 1691 27016 10060
rect 28482 10054 28602 10060
rect 30215 1882 30325 1886
rect 29682 1762 29688 1882
rect 29808 1877 30330 1882
rect 29808 1767 30215 1877
rect 30325 1767 30330 1877
rect 29808 1762 30330 1767
rect 30215 1758 30325 1762
rect 26892 1581 26901 1691
rect 27011 1581 27020 1691
rect 26896 1576 27016 1581
<< via2 >>
rect 28044 29470 28100 29526
rect 31367 29297 31657 29587
rect 26477 10675 26587 10785
rect 30215 1767 30325 1877
rect 26901 1581 27011 1691
<< metal3 >>
rect 3181 42932 3479 42937
rect 3180 42931 31662 42932
rect 3180 42633 3181 42931
rect 3479 42633 31662 42931
rect 3180 42632 31662 42633
rect 3181 42627 3479 42632
rect 28034 31298 28040 31362
rect 28104 31298 28110 31362
rect 28042 29531 28102 31298
rect 31362 29587 31662 42632
rect 28039 29526 28105 29531
rect 28039 29470 28044 29526
rect 28100 29470 28105 29526
rect 28039 29465 28105 29470
rect 31362 29297 31367 29587
rect 31657 29297 31662 29587
rect 31362 29292 31662 29297
rect 23981 10790 24099 10795
rect 23980 10789 26592 10790
rect 23980 10671 23981 10789
rect 24099 10785 26592 10789
rect 24099 10675 26477 10785
rect 26587 10675 26592 10785
rect 24099 10671 26592 10675
rect 23980 10670 26592 10671
rect 23981 10665 24099 10670
rect 30210 1877 31432 1882
rect 30210 1767 30215 1877
rect 30325 1767 31432 1877
rect 30210 1762 31432 1767
rect 26896 1691 27016 1696
rect 26896 1581 26901 1691
rect 27011 1581 27016 1691
rect 26896 1203 27016 1581
rect 31312 1343 31432 1762
rect 31307 1225 31313 1343
rect 31431 1225 31437 1343
rect 31312 1224 31432 1225
rect 26891 1085 26897 1203
rect 27015 1085 27021 1203
rect 26896 1084 27016 1085
<< via3 >>
rect 3181 42633 3479 42931
rect 28040 31298 28104 31362
rect 23981 10671 24099 10789
rect 31313 1225 31431 1343
rect 26897 1085 27015 1203
<< metal4 >>
rect 200 42932 500 44152
rect 798 43950 858 45152
rect 1534 43950 1594 45152
rect 2270 43950 2330 45152
rect 3006 43950 3066 45152
rect 3742 43950 3802 45152
rect 4478 43950 4538 45152
rect 5214 43950 5274 45152
rect 5950 43950 6010 45152
rect 6686 43950 6746 45152
rect 7422 43950 7482 45152
rect 8158 43950 8218 45152
rect 8894 43950 8954 45152
rect 9630 43950 9690 45152
rect 9800 43950 10100 44152
rect 798 43944 10100 43950
rect 10366 43944 10426 45152
rect 11102 43944 11162 45152
rect 11838 43944 11898 45152
rect 12574 43944 12634 45152
rect 13310 43944 13370 45152
rect 14046 43944 14106 45152
rect 14782 43944 14842 45152
rect 15518 43944 15578 45152
rect 16254 43944 16314 45152
rect 16990 43944 17050 45152
rect 17726 43944 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 798 43890 28102 43944
rect 9800 43884 28102 43890
rect 200 42931 3480 42932
rect 200 42633 3181 42931
rect 3479 42633 3480 42931
rect 200 42632 3480 42633
rect 200 1000 500 42632
rect 9800 1000 10100 43884
rect 28042 31363 28102 43884
rect 28039 31362 28105 31363
rect 28039 31298 28040 31362
rect 28104 31298 28105 31362
rect 28039 31297 28105 31298
rect 22480 10789 24100 10790
rect 22480 10671 23981 10789
rect 24099 10671 24100 10789
rect 22480 10670 24100 10671
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 10670
rect 31312 1343 31432 1344
rect 31312 1225 31313 1343
rect 31431 1225 31432 1343
rect 26896 1203 27016 1204
rect 26896 1085 26897 1203
rect 27015 1085 27016 1203
rect 26896 0 27016 1085
rect 31312 0 31432 1225
use p3_opamp  p3_opamp_0
timestamp 1712865377
transform 0 1 31042 -1 0 19722
box 1516 -3504 16136 620
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
