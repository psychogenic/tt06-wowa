* NGSPICE file created from onehot2mux.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_lvt_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_4QFWD3 a_n93_n200# a_n35_n297# a_35_n200# w_n231_n419#
X0 a_35_n200# a_n35_n297# a_n93_n200# w_n231_n419# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.35
**devattr s=23200,916 d=23200,916
.ends

.subckt lvtnot a y VCCPIN VSUBS
XXM1 VSUBS a y VSUBS sky130_fd_pr__nfet_01v8_lvt_648S5X
XXM2 VCCPIN a y VCCPIN sky130_fd_pr__pfet_01v8_lvt_4QFWD3
.ends

.subckt sky130_fd_pr__nfet_01v8_Q7AWK3 a_n180_n374# a_20_n200# a_n78_n200# a_n33_n288#
X0 a_20_n200# a_n33_n288# a_n78_n200# a_n180_n374# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
**devattr s=23200,916 d=23200,916
.ends

.subckt sky130_fd_pr__pfet_01v8_SKB8XJ w_n216_n419# a_n33_n297# a_20_n200# a_n78_n200#
X0 a_20_n200# a_n33_n297# a_n78_n200# w_n216_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.2
**devattr s=23200,916 d=23200,916
.ends

.subckt passgate A Z GP GN VCCBPIN VSUBS
XXM1 VSUBS Z A GN sky130_fd_pr__nfet_01v8_Q7AWK3
XXM2 VCCBPIN GP A Z sky130_fd_pr__pfet_01v8_SKB8XJ
.ends

.subckt onehot2mux SEL IN0 IN1 OUT VCC VSS
Xx1 SEL SEL_N VCC VSS lvtnot
Xx2 IN1 OUT SEL_N SEL VCC VSS passgate
Xx3 IN0 OUT SEL SEL_N VCC VSS passgate
.ends

