magic
tech sky130A
magscale 1 2
timestamp 1713160935
<< metal1 >>
rect -18980 -430 -16960 0
rect -13400 -30 -13200 0
rect -13400 -180 -13370 -30
rect -13220 -180 -13200 -30
rect -13400 -200 -13200 -180
rect -11400 -20 -11200 0
rect -11400 -180 -11380 -20
rect -11220 -180 -11200 -20
rect -11400 -200 -11200 -180
rect -17780 -2130 -17770 -1990
rect -17600 -2130 -17590 -1990
rect -16180 -3430 -16170 -3270
rect -16020 -3430 -16010 -3270
rect -15130 -3480 -15120 -3320
rect -14960 -3480 -14950 -3320
rect -10940 -4270 -10500 -4170
rect -11030 -4550 -11020 -4270
rect -19190 -4800 -18670 -4560
rect -19200 -5000 -18670 -4800
rect -11315 -4910 -11020 -4550
rect -10840 -4910 -10500 -4270
rect -11315 -4990 -10500 -4910
rect -11202 -5170 -10857 -5108
rect -11202 -5380 -11150 -5170
rect -10900 -5380 -10857 -5170
rect -19210 -6000 -11530 -5800
rect -19210 -6020 -17600 -6000
rect -18200 -6130 -18000 -6120
rect -18200 -6190 -18180 -6130
rect -18020 -6190 -18000 -6130
rect -17950 -6140 -17600 -6020
rect -15740 -6040 -11530 -6000
rect -19200 -6233 -19000 -6200
rect -18200 -6233 -18000 -6190
rect -19200 -6366 -17984 -6233
rect -19200 -6400 -19000 -6366
rect -18200 -6370 -18000 -6366
rect -18550 -6490 -17720 -6470
rect -19200 -6670 -17720 -6490
rect -12990 -6630 -12690 -6040
rect -12380 -6630 -12080 -6040
rect -11830 -6630 -11530 -6040
rect -11202 -5870 -10857 -5380
rect -11202 -5900 -10540 -5870
rect -19200 -6690 -18350 -6670
rect -19200 -6800 -19000 -6690
rect -19200 -7000 -18110 -6860
rect -19200 -7140 -18780 -7000
rect -18390 -7140 -18110 -7000
rect -19200 -7200 -18110 -7140
rect -11202 -6890 -11000 -5900
rect -10850 -6890 -10540 -5900
rect -11202 -6950 -10540 -6890
rect -12350 -7550 -12340 -7250
rect -12160 -7550 -12150 -7250
rect -11202 -7325 -10857 -6950
rect -11425 -7380 -10857 -7325
rect -11730 -7600 -10857 -7380
rect -19200 -7710 -18070 -7600
rect -11425 -7655 -10857 -7600
rect -11202 -7662 -10857 -7655
rect -19200 -7800 -17460 -7710
rect -19190 -7970 -17460 -7800
rect -18210 -8240 -17840 -7970
rect -17240 -8240 -16870 -7920
rect -16560 -8240 -16190 -7870
rect -11025 -8050 -10755 -8005
rect -18210 -8600 -13000 -8240
rect -11025 -8315 -11000 -8050
rect -11780 -8550 -11000 -8315
rect -10790 -8550 -10755 -8050
rect -11780 -8585 -10755 -8550
rect -11780 -8600 -11510 -8585
<< via1 >>
rect -13370 -180 -13220 -30
rect -11380 -180 -11220 -20
rect -17770 -2130 -17600 -1990
rect -16170 -3430 -16020 -3270
rect -15120 -3480 -14960 -3320
rect -11020 -4910 -10840 -4270
rect -11150 -5380 -10900 -5170
rect -18180 -6190 -18020 -6130
rect -18780 -7140 -18390 -7000
rect -11000 -6890 -10850 -5900
rect -12340 -7550 -12160 -7250
rect -11000 -8550 -10790 -8050
<< metal2 >>
rect -13390 -30 -13210 -10
rect -13390 -180 -13370 -30
rect -13220 -71 -13210 -30
rect -11400 -20 -11210 -10
rect -13220 -180 -13206 -71
rect -13390 -310 -13206 -180
rect -13380 -314 -13206 -310
rect -11400 -180 -11380 -20
rect -11220 -180 -11210 -20
rect -11400 -270 -11210 -180
rect -13380 -1030 -13210 -314
rect -11400 -380 -11390 -270
rect -11230 -380 -11210 -270
rect -11400 -400 -11210 -380
rect -18110 -1990 -17570 -1950
rect -18110 -2040 -17770 -1990
rect -18110 -2180 -18070 -2040
rect -17840 -2130 -17770 -2040
rect -17600 -2130 -17570 -1990
rect -17840 -2140 -17570 -2130
rect -17840 -2180 -17800 -2140
rect -18110 -2200 -17800 -2180
rect -11420 -2450 -11240 -2440
rect -11420 -2580 -11380 -2450
rect -11260 -2580 -11240 -2450
rect -11420 -2820 -11240 -2580
rect -16210 -3270 -15970 -3230
rect -16210 -3430 -16170 -3270
rect -16020 -3430 -15970 -3270
rect -16210 -3580 -15970 -3430
rect -16210 -3730 -16170 -3580
rect -16000 -3730 -15970 -3580
rect -15150 -3320 -14940 -3290
rect -15150 -3480 -15120 -3320
rect -14960 -3480 -14940 -3320
rect -15150 -3540 -14940 -3480
rect -15150 -3680 -15130 -3540
rect -14970 -3680 -14940 -3540
rect -15150 -3700 -14940 -3680
rect -16210 -3740 -15970 -3730
rect -14580 -3860 -14450 -3660
rect -11070 -4270 -10520 -4200
rect -18122 -4870 -17797 -4838
rect -18122 -5070 -18090 -4870
rect -17840 -5070 -17797 -4870
rect -11070 -4910 -11020 -4270
rect -10840 -4910 -10730 -4270
rect -10590 -4910 -10520 -4270
rect -11070 -4960 -10520 -4910
rect -18122 -5112 -17797 -5070
rect -11900 -5112 -10860 -5110
rect -18122 -5170 -10860 -5112
rect -18122 -5380 -11150 -5170
rect -10900 -5380 -10860 -5170
rect -18122 -5437 -10860 -5380
rect -11900 -5440 -10860 -5437
rect -18200 -5880 -18000 -5850
rect -18200 -6010 -18180 -5880
rect -18020 -6010 -18000 -5880
rect -18200 -6130 -18000 -6010
rect -18200 -6190 -18180 -6130
rect -18020 -6190 -18000 -6130
rect -18200 -6210 -18000 -6190
rect -11050 -5900 -10570 -5860
rect -18710 -6880 -18500 -6840
rect -18710 -6980 -18680 -6880
rect -18530 -6980 -18500 -6880
rect -11050 -6890 -11000 -5900
rect -10850 -5910 -10570 -5900
rect -10850 -6890 -10770 -5910
rect -11050 -6900 -10770 -6890
rect -10620 -6900 -10570 -5910
rect -11050 -6950 -10570 -6900
rect -18710 -6990 -18500 -6980
rect -18780 -7000 -18390 -6990
rect -18780 -7150 -18390 -7140
rect -12380 -7060 -12150 -7030
rect -12380 -7220 -12360 -7060
rect -12170 -7220 -12150 -7060
rect -12380 -7250 -12150 -7220
rect -12380 -7550 -12340 -7250
rect -12160 -7550 -12150 -7250
rect -12380 -7560 -12150 -7550
rect -13900 -7850 -13190 -7840
rect -13900 -8000 -13880 -7850
rect -13740 -8000 -13190 -7850
rect -13900 -8010 -13190 -8000
rect -11025 -8010 -10755 -8005
rect -11030 -8040 -10500 -8010
rect -11030 -8050 -10720 -8040
rect -11030 -8550 -11000 -8050
rect -10790 -8550 -10720 -8050
rect -11030 -8570 -10720 -8550
rect -10540 -8570 -10500 -8040
rect -11030 -8600 -10500 -8570
<< via2 >>
rect -11390 -380 -11230 -270
rect -18070 -2180 -17840 -2040
rect -11380 -2580 -11260 -2450
rect -16170 -3730 -16000 -3580
rect -15130 -3680 -14970 -3540
rect -18090 -5070 -17840 -4870
rect -10730 -4910 -10590 -4270
rect -18180 -6010 -18020 -5880
rect -18680 -6980 -18530 -6880
rect -10770 -6900 -10620 -5910
rect -12360 -7220 -12170 -7060
rect -13880 -8000 -13740 -7850
rect -10720 -8570 -10540 -8040
<< metal3 >>
rect -11400 -270 -11220 -260
rect -11400 -380 -11390 -270
rect -11230 -380 -11220 -270
rect -18120 -2040 -17800 -2000
rect -18120 -2180 -18070 -2040
rect -17840 -2078 -17800 -2040
rect -11400 -2074 -11220 -380
rect -17840 -2180 -17795 -2078
rect -18120 -4870 -17795 -2180
rect -11475 -2450 -11144 -2074
rect -11475 -2580 -11380 -2450
rect -11260 -2580 -11144 -2450
rect -15150 -3540 -14940 -3500
rect -18120 -5070 -18090 -4870
rect -17840 -5070 -17795 -4870
rect -18120 -5100 -17795 -5070
rect -16210 -3580 -15970 -3550
rect -16210 -3730 -16170 -3580
rect -16000 -3730 -15970 -3580
rect -18710 -5450 -17070 -5430
rect -18710 -5580 -18690 -5450
rect -18520 -5580 -17070 -5450
rect -16210 -5540 -15970 -3730
rect -15150 -3680 -15130 -3540
rect -14970 -3680 -14940 -3540
rect -15150 -3900 -14940 -3680
rect -15150 -4110 -14490 -3900
rect -18710 -5585 -17070 -5580
rect -16790 -5585 -15970 -5540
rect -18710 -5600 -15970 -5585
rect -18200 -5720 -18000 -5700
rect -18200 -5840 -18170 -5720
rect -18020 -5840 -18000 -5720
rect -17255 -5755 -15970 -5600
rect -16790 -5780 -15970 -5755
rect -18200 -5880 -18000 -5840
rect -18200 -6010 -18180 -5880
rect -18020 -6010 -18000 -5880
rect -18200 -6040 -18000 -6010
rect -18710 -6760 -18500 -6740
rect -18710 -6860 -18680 -6760
rect -18530 -6860 -18500 -6760
rect -18710 -6880 -18500 -6860
rect -18710 -6970 -18680 -6880
rect -18690 -6980 -18680 -6970
rect -18530 -6970 -18500 -6880
rect -18530 -6980 -18520 -6970
rect -18690 -6985 -18520 -6980
rect -14760 -7240 -14490 -4110
rect -13880 -5450 -13700 -5430
rect -13880 -5570 -13850 -5450
rect -13720 -5570 -13700 -5450
rect -13880 -5700 -13700 -5570
rect -13878 -7830 -13752 -5700
rect -11475 -6000 -11144 -2580
rect -10780 -4220 -10590 -4200
rect -10780 -4240 -10390 -4220
rect -10780 -4270 -9160 -4240
rect -10780 -4910 -10730 -4270
rect -10590 -4910 -9160 -4270
rect -10780 -4960 -9160 -4910
rect -10570 -4970 -9160 -4960
rect -10800 -5910 -10300 -5870
rect -12380 -6230 -11140 -6000
rect -12380 -7060 -12140 -6230
rect -10800 -6900 -10770 -5910
rect -10620 -5920 -10300 -5910
rect -10620 -6900 -10530 -5920
rect -10350 -6900 -10300 -5920
rect -10800 -6950 -10300 -6900
rect -12380 -7220 -12360 -7060
rect -12170 -7220 -12140 -7060
rect -12380 -7240 -12140 -7220
rect -13900 -7850 -13710 -7830
rect -13900 -8000 -13880 -7850
rect -13740 -8000 -13710 -7850
rect -13900 -8020 -13710 -8000
rect -11030 -8040 -9220 -8010
rect -11030 -8570 -10720 -8040
rect -10540 -8570 -9220 -8040
rect -11030 -8590 -9220 -8570
rect -10780 -8600 -9220 -8590
rect -10490 -8610 -9220 -8600
<< via3 >>
rect -18690 -5580 -18520 -5450
rect -18170 -5840 -18020 -5720
rect -18680 -6860 -18530 -6760
rect -13850 -5570 -13720 -5450
rect -10530 -6900 -10350 -5920
<< metal4 >>
rect -13879 -5274 -13701 -5251
rect -18166 -5407 -13701 -5274
rect -18710 -5450 -18500 -5410
rect -18710 -5580 -18690 -5450
rect -18520 -5580 -18500 -5450
rect -18166 -5480 -18033 -5407
rect -13879 -5450 -13701 -5407
rect -18710 -6760 -18500 -5580
rect -18200 -5720 -18000 -5480
rect -13879 -5570 -13850 -5450
rect -13720 -5570 -13701 -5450
rect -13879 -5599 -13701 -5570
rect -18200 -5840 -18170 -5720
rect -18020 -5840 -18000 -5720
rect -18200 -5850 -18000 -5840
rect -18710 -6860 -18680 -6760
rect -18530 -6860 -18500 -6760
rect -10810 -5880 -10320 -5870
rect -10810 -5920 -9650 -5880
rect -18681 -6861 -18529 -6860
rect -10810 -6900 -10530 -5920
rect -10350 -6900 -9650 -5920
rect -10810 -6920 -9650 -6900
rect -10810 -6950 -10320 -6920
use comparator_stefan  x1
timestamp 1713150544
transform 1 0 -28445 0 1 -10990
box 9445 5990 17870 10730
use analogswitch  x2
timestamp 1713149804
transform 1 0 -18620 0 1 -12120
box 5220 3520 7200 5620
use onehot2mux  x3
timestamp 1713137925
transform 1 0 -17650 0 1 -9780
box -550 1780 3445 3920
use sky130_fd_pr__cap_mim_m3_1_4HHTN9  XC1
timestamp 1713158458
transform 1 0 -8824 0 1 -4130
box -1186 -4640 1186 4640
<< labels >>
flabel metal1 -19200 -5000 -19000 -4800 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
flabel metal1 -18600 -200 -18400 0 0 FreeSans 1280 0 0 0 VCC
port 0 nsew
flabel metal1 -13400 -200 -13200 0 0 FreeSans 1280 0 0 0 EN_N
port 6 nsew
flabel metal1 -11400 -200 -11200 0 0 FreeSans 1280 0 0 0 RESULT
port 5 nsew
flabel metal1 -19200 -7200 -19000 -7000 0 FreeSans 1280 0 0 0 THRESHV
port 3 nsew
flabel metal1 -19200 -6800 -19000 -6600 0 FreeSans 1280 0 0 0 INPUT
port 2 nsew
flabel metal1 -19200 -6400 -19000 -6200 0 FreeSans 1280 0 0 0 CALIB
port 4 nsew
flabel metal1 -19200 -6000 -19000 -5800 0 FreeSans 1280 0 0 0 VCC
port 0 nsew
flabel metal1 -19200 -7800 -19000 -7600 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
<< end >>
