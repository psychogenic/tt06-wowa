magic
tech sky130A
magscale 1 2
timestamp 1713118242
<< error_s >>
rect 369 10666 422 10667
rect 1160 10666 1213 10667
rect 351 10632 422 10666
rect 1142 10632 1213 10666
rect 352 10631 422 10632
rect 1143 10631 1213 10632
rect 369 10597 440 10631
rect 1160 10597 1231 10631
rect 182 10564 240 10570
rect 182 10530 194 10564
rect 182 10524 240 10530
rect 182 10370 240 10376
rect 182 10336 194 10370
rect 182 10330 240 10336
rect 369 10234 439 10597
rect 973 10564 1031 10570
rect 551 10529 609 10535
rect 973 10530 985 10564
rect 551 10495 563 10529
rect 973 10524 1031 10530
rect 551 10489 609 10495
rect 973 10370 1031 10376
rect 973 10336 985 10370
rect 973 10330 1031 10336
rect 551 10317 609 10323
rect 551 10283 563 10317
rect 551 10277 609 10283
rect 1160 10234 1230 10597
rect 1342 10529 1400 10535
rect 1342 10495 1354 10529
rect 1342 10489 1400 10495
rect 1342 10317 1400 10323
rect 1342 10283 1354 10317
rect 1342 10277 1400 10283
rect 369 10198 422 10234
rect 1160 10198 1213 10234
rect 1973 5999 2008 6016
rect 1974 5998 2008 5999
rect 1974 5962 2044 5998
rect 1782 5931 1844 5937
rect 1782 5897 1794 5931
rect 1991 5928 2062 5962
rect 1782 5891 1844 5897
rect 1782 5719 1844 5725
rect 1414 5616 1582 5715
rect 1782 5685 1794 5719
rect 1782 5679 1844 5685
rect 369 5615 422 5616
rect 1160 5615 1213 5616
rect 351 5581 422 5615
rect 1142 5581 1213 5615
rect 352 5580 422 5581
rect 1143 5580 1213 5581
rect 1991 5583 2061 5928
rect 2173 5860 2231 5866
rect 2173 5826 2185 5860
rect 2173 5820 2231 5826
rect 2173 5666 2231 5672
rect 2173 5632 2185 5666
rect 2173 5626 2231 5632
rect 369 5546 440 5580
rect 1160 5546 1231 5580
rect 1991 5547 2044 5583
rect 182 5513 240 5519
rect 182 5479 194 5513
rect 182 5473 240 5479
rect 182 5319 240 5325
rect 182 5285 194 5319
rect 182 5279 240 5285
rect 369 5183 439 5546
rect 973 5513 1031 5519
rect 551 5478 609 5484
rect 973 5479 985 5513
rect 551 5444 563 5478
rect 973 5473 1031 5479
rect 551 5438 609 5444
rect 973 5319 1031 5325
rect 973 5285 985 5319
rect 973 5279 1031 5285
rect 551 5266 609 5272
rect 551 5232 563 5266
rect 551 5226 609 5232
rect 1160 5183 1230 5546
rect 1342 5478 1400 5484
rect 1342 5444 1354 5478
rect 1342 5438 1400 5444
rect 1342 5266 1400 5272
rect 1342 5232 1354 5266
rect 1342 5226 1400 5232
rect 369 5147 422 5183
rect 1160 5147 1213 5183
use passgate  x1
array 0 0 791 0 1 5051
timestamp 1713118242
transform 1 0 53 0 1 4600
box -53 -4000 738 1051
use passgate  x3
array 0 0 791 0 1 5051
timestamp 1713118242
transform 1 0 844 0 1 4600
box -53 -4000 738 1051
use lvtnot  x5
timestamp 1713118242
transform 1 0 1635 0 1 5000
box -53 -4400 778 1069
<< end >>
