magic
tech sky130A
timestamp 1712893257
<< pwell >>
rect -885 -155 885 155
<< nmos >>
rect -787 -50 -587 50
rect -558 -50 -358 50
rect -329 -50 -129 50
rect -100 -50 100 50
rect 129 -50 329 50
rect 358 -50 558 50
rect 587 -50 787 50
<< ndiff >>
rect -816 44 -787 50
rect -816 -44 -810 44
rect -793 -44 -787 44
rect -816 -50 -787 -44
rect -587 44 -558 50
rect -587 -44 -581 44
rect -564 -44 -558 44
rect -587 -50 -558 -44
rect -358 44 -329 50
rect -358 -44 -352 44
rect -335 -44 -329 44
rect -358 -50 -329 -44
rect -129 44 -100 50
rect -129 -44 -123 44
rect -106 -44 -100 44
rect -129 -50 -100 -44
rect 100 44 129 50
rect 100 -44 106 44
rect 123 -44 129 44
rect 100 -50 129 -44
rect 329 44 358 50
rect 329 -44 335 44
rect 352 -44 358 44
rect 329 -50 358 -44
rect 558 44 587 50
rect 558 -44 564 44
rect 581 -44 587 44
rect 558 -50 587 -44
rect 787 44 816 50
rect 787 -44 793 44
rect 810 -44 816 44
rect 787 -50 816 -44
<< ndiffc >>
rect -810 -44 -793 44
rect -581 -44 -564 44
rect -352 -44 -335 44
rect -123 -44 -106 44
rect 106 -44 123 44
rect 335 -44 352 44
rect 564 -44 581 44
rect 793 -44 810 44
<< psubdiff >>
rect -867 120 -819 137
rect 819 120 867 137
rect -867 89 -850 120
rect 850 89 867 120
rect -867 -120 -850 -89
rect 850 -120 867 -89
rect -867 -137 -819 -120
rect 819 -137 867 -120
<< psubdiffcont >>
rect -819 120 819 137
rect -867 -89 -850 89
rect 850 -89 867 89
rect -819 -137 819 -120
<< poly >>
rect -787 86 -587 94
rect -787 69 -779 86
rect -595 69 -587 86
rect -787 50 -587 69
rect -558 86 -358 94
rect -558 69 -550 86
rect -366 69 -358 86
rect -558 50 -358 69
rect -329 86 -129 94
rect -329 69 -321 86
rect -137 69 -129 86
rect -329 50 -129 69
rect -100 86 100 94
rect -100 69 -92 86
rect 92 69 100 86
rect -100 50 100 69
rect 129 86 329 94
rect 129 69 137 86
rect 321 69 329 86
rect 129 50 329 69
rect 358 86 558 94
rect 358 69 366 86
rect 550 69 558 86
rect 358 50 558 69
rect 587 86 787 94
rect 587 69 595 86
rect 779 69 787 86
rect 587 50 787 69
rect -787 -69 -587 -50
rect -787 -86 -779 -69
rect -595 -86 -587 -69
rect -787 -94 -587 -86
rect -558 -69 -358 -50
rect -558 -86 -550 -69
rect -366 -86 -358 -69
rect -558 -94 -358 -86
rect -329 -69 -129 -50
rect -329 -86 -321 -69
rect -137 -86 -129 -69
rect -329 -94 -129 -86
rect -100 -69 100 -50
rect -100 -86 -92 -69
rect 92 -86 100 -69
rect -100 -94 100 -86
rect 129 -69 329 -50
rect 129 -86 137 -69
rect 321 -86 329 -69
rect 129 -94 329 -86
rect 358 -69 558 -50
rect 358 -86 366 -69
rect 550 -86 558 -69
rect 358 -94 558 -86
rect 587 -69 787 -50
rect 587 -86 595 -69
rect 779 -86 787 -69
rect 587 -94 787 -86
<< polycont >>
rect -779 69 -595 86
rect -550 69 -366 86
rect -321 69 -137 86
rect -92 69 92 86
rect 137 69 321 86
rect 366 69 550 86
rect 595 69 779 86
rect -779 -86 -595 -69
rect -550 -86 -366 -69
rect -321 -86 -137 -69
rect -92 -86 92 -69
rect 137 -86 321 -69
rect 366 -86 550 -69
rect 595 -86 779 -69
<< locali >>
rect -867 120 -819 137
rect 819 120 867 137
rect -867 89 -850 120
rect 850 89 867 120
rect -787 69 -779 86
rect -595 69 -587 86
rect -558 69 -550 86
rect -366 69 -358 86
rect -329 69 -321 86
rect -137 69 -129 86
rect -100 69 -92 86
rect 92 69 100 86
rect 129 69 137 86
rect 321 69 329 86
rect 358 69 366 86
rect 550 69 558 86
rect 587 69 595 86
rect 779 69 787 86
rect -810 44 -793 52
rect -810 -52 -793 -44
rect -581 44 -564 52
rect -581 -52 -564 -44
rect -352 44 -335 52
rect -352 -52 -335 -44
rect -123 44 -106 52
rect -123 -52 -106 -44
rect 106 44 123 52
rect 106 -52 123 -44
rect 335 44 352 52
rect 335 -52 352 -44
rect 564 44 581 52
rect 564 -52 581 -44
rect 793 44 810 52
rect 793 -52 810 -44
rect -787 -86 -779 -69
rect -595 -86 -587 -69
rect -558 -86 -550 -69
rect -366 -86 -358 -69
rect -329 -86 -321 -69
rect -137 -86 -129 -69
rect -100 -86 -92 -69
rect 92 -86 100 -69
rect 129 -86 137 -69
rect 321 -86 329 -69
rect 358 -86 366 -69
rect 550 -86 558 -69
rect 587 -86 595 -69
rect 779 -86 787 -69
rect -867 -120 -850 -89
rect 850 -120 867 -89
rect -867 -137 -819 -120
rect 819 -137 867 -120
<< viali >>
rect -779 69 -595 86
rect -550 69 -366 86
rect -321 69 -137 86
rect -92 69 92 86
rect 137 69 321 86
rect 366 69 550 86
rect 595 69 779 86
rect -810 -44 -793 44
rect -581 -44 -564 44
rect -352 -44 -335 44
rect -123 -44 -106 44
rect 106 -44 123 44
rect 335 -44 352 44
rect 564 -44 581 44
rect 793 -44 810 44
rect -779 -86 -595 -69
rect -550 -86 -366 -69
rect -321 -86 -137 -69
rect -92 -86 92 -69
rect 137 -86 321 -69
rect 366 -86 550 -69
rect 595 -86 779 -69
<< metal1 >>
rect -785 86 -589 89
rect -785 69 -779 86
rect -595 69 -589 86
rect -785 66 -589 69
rect -556 86 -360 89
rect -556 69 -550 86
rect -366 69 -360 86
rect -556 66 -360 69
rect -327 86 -131 89
rect -327 69 -321 86
rect -137 69 -131 86
rect -327 66 -131 69
rect -98 86 98 89
rect -98 69 -92 86
rect 92 69 98 86
rect -98 66 98 69
rect 131 86 327 89
rect 131 69 137 86
rect 321 69 327 86
rect 131 66 327 69
rect 360 86 556 89
rect 360 69 366 86
rect 550 69 556 86
rect 360 66 556 69
rect 589 86 785 89
rect 589 69 595 86
rect 779 69 785 86
rect 589 66 785 69
rect -813 44 -790 50
rect -813 -44 -810 44
rect -793 -44 -790 44
rect -813 -50 -790 -44
rect -584 44 -561 50
rect -584 -44 -581 44
rect -564 -44 -561 44
rect -584 -50 -561 -44
rect -355 44 -332 50
rect -355 -44 -352 44
rect -335 -44 -332 44
rect -355 -50 -332 -44
rect -126 44 -103 50
rect -126 -44 -123 44
rect -106 -44 -103 44
rect -126 -50 -103 -44
rect 103 44 126 50
rect 103 -44 106 44
rect 123 -44 126 44
rect 103 -50 126 -44
rect 332 44 355 50
rect 332 -44 335 44
rect 352 -44 355 44
rect 332 -50 355 -44
rect 561 44 584 50
rect 561 -44 564 44
rect 581 -44 584 44
rect 561 -50 584 -44
rect 790 44 813 50
rect 790 -44 793 44
rect 810 -44 813 44
rect 790 -50 813 -44
rect -785 -69 -589 -66
rect -785 -86 -779 -69
rect -595 -86 -589 -69
rect -785 -89 -589 -86
rect -556 -69 -360 -66
rect -556 -86 -550 -69
rect -366 -86 -360 -69
rect -556 -89 -360 -86
rect -327 -69 -131 -66
rect -327 -86 -321 -69
rect -137 -86 -131 -69
rect -327 -89 -131 -86
rect -98 -69 98 -66
rect -98 -86 -92 -69
rect 92 -86 98 -69
rect -98 -89 98 -86
rect 131 -69 327 -66
rect 131 -86 137 -69
rect 321 -86 327 -69
rect 131 -89 327 -86
rect 360 -69 556 -66
rect 360 -86 366 -69
rect 550 -86 556 -69
rect 360 -89 556 -86
rect 589 -69 785 -66
rect 589 -86 595 -69
rect 779 -86 785 -69
rect 589 -89 785 -86
<< properties >>
string FIXED_BBOX -858 -128 858 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 2.0 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
